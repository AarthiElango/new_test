module adder(a,b,c); //DUT code start
input [15:0] a,b;
output [16:0] c;

assign c = a + b;

endmodule //DUT code end